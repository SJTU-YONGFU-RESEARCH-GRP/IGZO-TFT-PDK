VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO INV_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN INV_1 0 -0.15 ;
  SIZE 4.5 BY 5.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.05 1.8 1.35 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 2.85 4.2 3.15 ;
        RECT 2.7 1.65 4.2 1.95 ;
        RECT 3.3 1.65 3.6 3.15 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 4.65 4.5 4.95 ;
        RECT 0.3 4.05 4.2 4.35 ;
        RECT 2.1 4.05 2.4 4.95 ;
        RECT 0.3 3.45 0.6 4.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 4.5 0.15 ;
        RECT 0.3 0.45 4.2 0.75 ;
        RECT 2.1 -0.15 2.4 0.75 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.1 3.45 3 3.75 ;
      RECT 2.1 2.85 2.4 3.75 ;
      RECT 0.3 2.85 2.4 3.15 ;
      RECT 0.9 1.65 1.2 3.15 ;
      RECT 0.3 1.65 1.8 1.95 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END INV_1

MACRO NAND2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN NAND2_1 0 -0.15 ;
  SIZE 7.6 BY 5.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.05 1.8 1.35 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 1.05 4.2 1.35 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 2.85 6.6 3.15 ;
        RECT 5.1 1.65 6.6 1.95 ;
        RECT 5.7 1.65 6 3.15 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 4.65 7.6 4.95 ;
        RECT 0.3 4.05 4.2 4.35 ;
        RECT 2.1 4.05 2.4 4.95 ;
        RECT 0.3 3.45 0.6 4.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 7.6 0.15 ;
        RECT 5.1 4.05 7.3 4.35 ;
        RECT 7 0.45 7.3 4.35 ;
        RECT 2.7 0.45 7.3 0.75 ;
        RECT 3.9 -0.15 4.2 0.75 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.1 1.65 4.2 1.95 ;
      RECT 2.1 0.45 2.4 1.95 ;
      RECT 0.3 0.45 2.4 0.75 ;
      RECT 2.1 3.45 3 3.75 ;
      RECT 2.1 2.85 2.4 3.75 ;
      RECT 0.3 2.85 2.4 3.15 ;
      RECT 0.9 1.65 1.2 3.15 ;
      RECT 0.3 1.65 1.8 1.95 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END NAND2_1

MACRO NOR2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN NOR2_1 0 -0.15 ;
  SIZE 7.5 BY 5.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 0.3 1.05 1.8 1.35 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 1.05 4.2 1.35 ;
    END
  END B
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 2.7 2.85 6.6 3.15 ;
        RECT 5.1 1.65 6.6 1.95 ;
        RECT 5.7 1.65 6 3.15 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 4.65 7.5 4.95 ;
        RECT 0.3 4.05 4.2 4.35 ;
        RECT 2.1 4.05 2.4 4.95 ;
        RECT 0.3 3.45 0.6 4.35 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 7.5 0.15 ;
        RECT 5.1 4.05 7.2 4.35 ;
        RECT 6.9 0.45 7.2 4.35 ;
        RECT 0.3 0.45 7.2 0.75 ;
        RECT 3.9 -0.15 4.2 0.75 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 2.1 3.45 3 3.75 ;
      RECT 2.1 2.85 2.4 3.75 ;
      RECT 0.3 2.85 2.4 3.15 ;
      RECT 0.9 1.65 1.2 3.15 ;
      RECT 0.3 1.65 4.2 1.95 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END NOR2_1

MACRO all
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN all 0 -0.15 ;
  SIZE 12.3 BY 11.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CTRL0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 7.65 2.1 7.95 ;
      LAYER Metal2 ;
        RECT 1.8 7.65 3 7.95 ;
        RECT 1.8 7.05 2.1 7.95 ;
      LAYER VIA1 ;
        RECT 1.85 7.7 2.05 7.9 ;
    END
  END CTRL0
  PIN CTRL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.8 9.45 8.7 9.75 ;
        RECT 8.4 8.55 8.7 9.75 ;
      LAYER VIA1 ;
        RECT 8.45 9.5 8.65 9.7 ;
    END
  END CTRL1
  PIN CTRL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.2 2.85 10.5 3.15 ;
      LAYER Metal2 ;
        RECT 10.2 2.85 10.5 3.75 ;
        RECT 9.3 2.85 10.5 3.15 ;
      LAYER VIA1 ;
        RECT 10.25 2.9 10.45 3.1 ;
    END
  END CTRL2
  PIN CTRL3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.6 1.05 4.5 1.35 ;
        RECT 3.6 1.05 3.9 2.25 ;
      LAYER VIA1 ;
        RECT 3.65 1.1 3.85 1.3 ;
    END
  END CTRL3
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.4 5.25 6.9 5.55 ;
        RECT 6 4.65 6.3 6.15 ;
      LAYER Metal2 ;
        RECT 5.4 5.25 6.9 5.55 ;
        RECT 6 4.65 6.3 6.15 ;
      LAYER VIA1 ;
        RECT 5.55 5.3 5.75 5.5 ;
        RECT 6.05 5.3 6.25 5.5 ;
        RECT 6.55 5.3 6.75 5.5 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 5.85 9.3 7.35 ;
        RECT 7.8 6.45 9.3 6.75 ;
        RECT 7.8 5.85 8.1 7.35 ;
        RECT 6.6 3.45 8.1 3.75 ;
        RECT 6.6 2.25 8.1 2.55 ;
        RECT 7.2 2.25 7.5 3.75 ;
        RECT 4.2 8.25 5.7 8.55 ;
        RECT 4.2 7.05 5.7 7.35 ;
        RECT 4.8 7.05 5.1 8.55 ;
        RECT 4.2 3.45 4.5 4.95 ;
        RECT 3 4.05 4.5 4.35 ;
        RECT 3 3.45 3.3 4.95 ;
      LAYER Metal2 ;
        RECT 3.6 7.65 8.7 7.95 ;
        RECT 8.4 6.45 8.7 7.95 ;
        RECT 3.6 2.85 7.5 3.15 ;
        RECT 3.6 2.85 3.9 7.95 ;
      LAYER VIA1 ;
        RECT 3.65 4.1 3.85 4.3 ;
        RECT 4.85 7.7 5.05 7.9 ;
        RECT 7.25 2.9 7.45 3.1 ;
        RECT 8.45 6.5 8.65 6.7 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 10.65 12.3 10.95 ;
        RECT 11.4 0.45 11.7 10.95 ;
        RECT 1.2 0.45 11.7 0.75 ;
        RECT 1.2 0.45 1.5 9.75 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 12.3 0.15 ;
        RECT 0.6 10.05 11.1 10.35 ;
        RECT 10.8 1.05 11.1 10.35 ;
        RECT 0.6 -0.15 0.9 10.35 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 10.2 1.05 10.5 1.95 ;
      RECT 6.6 1.05 10.5 1.35 ;
      RECT 9 3.45 10.5 3.75 ;
      RECT 9.6 2.25 9.9 3.75 ;
      RECT 8.4 2.25 10.5 2.55 ;
      RECT 8.4 1.65 8.7 2.55 ;
      RECT 7.8 1.65 8.7 1.95 ;
      RECT 9.6 9.45 10.5 9.75 ;
      RECT 10.2 5.85 10.5 9.75 ;
      RECT 9 7.65 9.3 9.75 ;
      RECT 7.8 8.25 8.1 9.75 ;
      RECT 7.8 8.85 9.3 9.15 ;
      RECT 9 7.65 9.9 7.95 ;
      RECT 9.6 7.05 9.9 7.95 ;
      RECT 1.8 9.45 5.7 9.75 ;
      RECT 1.8 8.85 2.1 9.75 ;
      RECT 2.4 2.85 2.7 3.75 ;
      RECT 2.4 2.85 3.3 3.15 ;
      RECT 3 1.05 3.3 3.15 ;
      RECT 4.2 1.05 4.5 2.55 ;
      RECT 3 1.65 4.5 1.95 ;
      RECT 3.6 8.85 4.5 9.15 ;
      RECT 3.6 8.25 3.9 9.15 ;
      RECT 1.8 8.25 3.9 8.55 ;
      RECT 2.4 7.05 2.7 8.55 ;
      RECT 1.8 7.05 3.3 7.35 ;
      RECT 1.8 1.05 2.1 4.95 ;
      RECT 1.8 1.05 2.7 1.35 ;
      RECT 6.6 4.65 10.5 4.95 ;
      RECT 6.6 5.85 6.9 9.75 ;
      RECT 5.4 1.05 5.7 4.95 ;
      RECT 1.8 5.85 5.7 6.15 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END all

END LIBRARY
