VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MANUFACTURINGGRID 0.005 ;

LAYER TopGate
  TYPE MASTERSLICE ;
END TopGate

LAYER BtmGate
  TYPE MASTERSLICE ;
END BtmGate

LAYER AA
  TYPE MASTERSLICE ;
END AA

LAYER Cont
  TYPE CUT ;
  SPACING 0.2 ;
  WIDTH 0.2 ;
END Cont

LAYER Metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  SPACING 0.3 ;
END Metal1

LAYER VIA1
  TYPE CUT ;
  SPACING 0.3 ;
  WIDTH 0.2 ;
END VIA1

LAYER Metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  SPACING 0.3 ;
END Metal2

LAYER VIA2
  TYPE CUT ;
  SPACING 0.3 ;
  WIDTH 0.2 ;
END VIA2

LAYER Metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  SPACING 0.3 ;
END Metal3

LAYER VIA3
  TYPE CUT ;
  SPACING 0.3 ;
  WIDTH 0.2 ;
END VIA3

LAYER Metal4
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  SPACING 0.3 ;
END Metal4

LAYER VIA4
  TYPE CUT ;
  SPACING 0.3 ;
  WIDTH 0.2 ;
END VIA4

LAYER Metal5
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  SPACING 0.3 ;
END Metal5

LAYER VIA5
  TYPE CUT ;
  SPACING 0.3 ;
  WIDTH 0.2 ;
END VIA5

LAYER Metal6
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 0.6 0.6 ;
  WIDTH 0.3 ;
  OFFSET 0.3 0.3 ;
  SPACING 0.3 ;
END Metal6

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA M6_M5 DEFAULT
  LAYER Metal5 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal6 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER VIA5 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    RESISTANCE 6.400000 ;
END M6_M5

VIA M5_M4 DEFAULT
  LAYER Metal4 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal5 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER VIA4 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    RESISTANCE 6.400000 ;
END M5_M4

VIA M4_M3  DEFAULT
  LAYER Metal3 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal4 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER VIA3 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    RESISTANCE 6.400000 ;
END M4_M3

VIA M3_M2  DEFAULT
  LAYER Metal2 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal3 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER VIA2 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    RESISTANCE 6.400000 ;
END M3_M2

VIA M2_M1  DEFAULT
  LAYER Metal1 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal2 ;
   RECT -0.15 -0.15 0.15 0.15 ;
  LAYER VIA1 ;
    RECT -0.1 -0.1 0.1 0.1 ;
    RESISTANCE 6.400000 ;
END M2_M1

VIA M1_TopGate 
  LAYER TopGate ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal1 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Cont ;
    RECT -0.1 -0.1 0.1 0.1 ;
END M1_TopGate

VIA M1_BtmGate 
  LAYER BtmGate ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal1 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Cont ;
    RECT -0.1 -0.1 0.1 0.1 ;
END M1_BtmGate

VIA M1_AA 
  LAYER AA ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Metal1 ;
    RECT -0.15 -0.15 0.15 0.15 ;
  LAYER Cont ;
    RECT -0.1 -0.1 0.1 0.1 ;
END M1_AA

SITE CoreSite
  CLASS CORE ;
  SIZE 0.6 BY 11.1 ;
END CoreSite

END LIBRARY
