VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO CatenaDesignType STRING ;
END PROPERTYDEFINITIONS

MACRO INV_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN INV_1 0 -0.15 ;
  SIZE 12.3 BY 11.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN CTRL0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 1.8 7.65 2.1 7.95 ;
      LAYER Metal2 ;
        RECT 1.8 7.65 3 7.95 ;
        RECT 1.8 7.05 2.1 7.95 ;
      LAYER VIA1 ;
        RECT 1.85 7.7 2.05 7.9 ;
    END
  END CTRL0
  PIN CTRL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 7.8 9.45 8.7 9.75 ;
        RECT 8.4 8.55 8.7 9.75 ;
      LAYER VIA1 ;
        RECT 8.45 9.5 8.65 9.7 ;
    END
  END CTRL1
  PIN CTRL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.2 2.85 10.5 3.15 ;
      LAYER Metal2 ;
        RECT 10.2 2.85 10.5 3.75 ;
        RECT 9.3 2.85 10.5 3.15 ;
      LAYER VIA1 ;
        RECT 10.25 2.9 10.45 3.1 ;
    END
  END CTRL2
  PIN CTRL3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 3.6 1.05 4.5 1.35 ;
        RECT 3.6 1.05 3.9 2.25 ;
      LAYER VIA1 ;
        RECT 3.65 1.1 3.85 1.3 ;
    END
  END CTRL3
  PIN IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 5.4 5.25 6.9 5.55 ;
        RECT 6 4.65 6.3 6.15 ;
      LAYER Metal2 ;
        RECT 5.4 5.25 6.9 5.55 ;
        RECT 6 4.65 6.3 6.15 ;
      LAYER VIA1 ;
        RECT 5.55 5.3 5.75 5.5 ;
        RECT 6.05 5.3 6.25 5.5 ;
        RECT 6.55 5.3 6.75 5.5 ;
    END
  END IN
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 5.85 9.3 7.35 ;
        RECT 7.8 6.45 9.3 6.75 ;
        RECT 7.8 5.85 8.1 7.35 ;
        RECT 6.6 3.45 8.1 3.75 ;
        RECT 6.6 2.25 8.1 2.55 ;
        RECT 7.2 2.25 7.5 3.75 ;
        RECT 4.2 8.25 5.7 8.55 ;
        RECT 4.2 7.05 5.7 7.35 ;
        RECT 4.8 7.05 5.1 8.55 ;
        RECT 4.2 3.45 4.5 4.95 ;
        RECT 3 4.05 4.5 4.35 ;
        RECT 3 3.45 3.3 4.95 ;
      LAYER Metal2 ;
        RECT 3.6 7.65 8.7 7.95 ;
        RECT 8.4 6.45 8.7 7.95 ;
        RECT 3.6 2.85 7.5 3.15 ;
        RECT 3.6 2.85 3.9 7.95 ;
      LAYER VIA1 ;
        RECT 3.65 4.1 3.85 4.3 ;
        RECT 4.85 7.7 5.05 7.9 ;
        RECT 7.25 2.9 7.45 3.1 ;
        RECT 8.45 6.5 8.65 6.7 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 10.65 12.3 10.95 ;
        RECT 11.4 0.45 11.7 10.95 ;
        RECT 1.2 0.45 11.7 0.75 ;
        RECT 1.2 0.45 1.5 9.75 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 12.3 0.15 ;
        RECT 0.6 10.05 11.1 10.35 ;
        RECT 10.8 1.05 11.1 10.35 ;
        RECT 0.6 -0.15 0.9 10.35 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 10.2 1.05 10.5 1.95 ;
      RECT 6.6 1.05 10.5 1.35 ;
      RECT 9 3.45 10.5 3.75 ;
      RECT 9.6 2.25 9.9 3.75 ;
      RECT 8.4 2.25 10.5 2.55 ;
      RECT 8.4 1.65 8.7 2.55 ;
      RECT 7.8 1.65 8.7 1.95 ;
      RECT 9.6 9.45 10.5 9.75 ;
      RECT 10.2 5.85 10.5 9.75 ;
      RECT 9 7.65 9.3 9.75 ;
      RECT 7.8 8.25 8.1 9.75 ;
      RECT 7.8 8.85 9.3 9.15 ;
      RECT 9 7.65 9.9 7.95 ;
      RECT 9.6 7.05 9.9 7.95 ;
      RECT 1.8 9.45 5.7 9.75 ;
      RECT 1.8 8.85 2.1 9.75 ;
      RECT 2.4 2.85 2.7 3.75 ;
      RECT 2.4 2.85 3.3 3.15 ;
      RECT 3 1.05 3.3 3.15 ;
      RECT 4.2 1.05 4.5 2.55 ;
      RECT 3 1.65 4.5 1.95 ;
      RECT 3.6 8.85 4.5 9.15 ;
      RECT 3.6 8.25 3.9 9.15 ;
      RECT 1.8 8.25 3.9 8.55 ;
      RECT 2.4 7.05 2.7 8.55 ;
      RECT 1.8 7.05 3.3 7.35 ;
      RECT 1.8 1.05 2.1 4.95 ;
      RECT 1.8 1.05 2.7 1.35 ;
      RECT 6.6 4.65 10.5 4.95 ;
      RECT 6.6 5.85 6.9 9.75 ;
      RECT 5.4 1.05 5.7 4.95 ;
      RECT 1.8 5.85 5.7 6.15 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END INV_1

MACRO NAND2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN NAND2_1 0 -0.15 ;
  SIZE 18.5 BY 11.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.1 5.25 9.4 6.155 ;
      LAYER Metal2 ;
        RECT 6.7 5.55 11.895 5.85 ;
        RECT 6.7 5.55 7 6.45 ;
      LAYER VIA1 ;
        RECT 9.15 5.6 9.35 5.8 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 13.4 5.25 14.2 5.55 ;
        RECT 4.3 5.25 5.1 5.55 ;
      LAYER Metal2 ;
        RECT 13.4 5.25 14.2 5.55 ;
        RECT 4.8 4.95 13.7 5.25 ;
        RECT 4.3 5.25 5.1 5.55 ;
      LAYER VIA1 ;
        RECT 4.85 5.3 5.05 5.5 ;
        RECT 13.45 5.3 13.65 5.5 ;
    END
  END B
  PIN CTRL0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 7.3 7.65 7.6 7.95 ;
      LAYER Metal2 ;
        RECT 7.3 7.65 8.2 7.95 ;
        RECT 7.3 7.35 7.6 7.95 ;
      LAYER VIA1 ;
        RECT 7.35 7.7 7.55 7.9 ;
    END
  END CTRL0
  PIN CTRL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 12.2 7.05 12.5 7.35 ;
      LAYER Metal2 ;
        RECT 11.9 7.05 12.8 7.35 ;
        RECT 12.5 6.75 12.8 7.35 ;
      LAYER VIA1 ;
        RECT 12.25 7.1 12.45 7.3 ;
    END
  END CTRL1
  PIN CTRL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 10.9 2.85 11.2 3.15 ;
      LAYER Metal2 ;
        RECT 10.9 2.85 11.8 3.15 ;
        RECT 10.9 2.85 11.2 3.45 ;
      LAYER VIA1 ;
        RECT 10.95 2.9 11.15 3.1 ;
    END
  END CTRL2
  PIN CTRL3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 3.6 2.85 3.9 3.15 ;
      LAYER Metal2 ;
        RECT 3.6 3.15 4.2 3.45 ;
        RECT 3.6 2.85 3.9 3.75 ;
      LAYER VIA1 ;
        RECT 3.65 2.9 3.85 3.1 ;
    END
  END CTRL3
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 14.5 3.45 16 3.75 ;
        RECT 12.1 2.25 16 2.55 ;
        RECT 15.1 2.25 15.4 3.75 ;
        RECT 15.2 8.25 15.5 9.75 ;
        RECT 14 8.85 15.5 9.15 ;
        RECT 14 7.65 14.3 9.75 ;
        RECT 10.4 7.65 14.3 7.95 ;
        RECT 10.4 7.65 10.7 9.75 ;
        RECT 4.2 2.85 8.1 3.15 ;
        RECT 7.8 1.05 8.1 3.15 ;
        RECT 4.2 1.05 4.5 3.15 ;
        RECT 3 1.65 4.5 1.95 ;
        RECT 3 1.05 3.3 2.55 ;
        RECT 2.5 8.25 6.4 8.55 ;
        RECT 2.5 7.05 4 7.35 ;
        RECT 3.1 7.05 3.4 8.55 ;
      LAYER Metal2 ;
        RECT 14.6 2.25 14.9 9.275 ;
        RECT 4 8.25 14.9 8.55 ;
        RECT 3.6 2.25 14.9 2.55 ;
        RECT 3.6 1.65 3.9 2.55 ;
      LAYER VIA1 ;
        RECT 3.65 1.7 3.85 1.9 ;
        RECT 4.35 8.3 4.55 8.5 ;
        RECT 13.95 2.3 14.15 2.5 ;
        RECT 14.65 8.9 14.85 9.1 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 10.65 18.5 10.95 ;
        RECT 17 0.45 17.3 9.75 ;
        RECT 0.6 0.45 17.3 0.75 ;
        RECT 9.7 1.05 13.6 1.35 ;
        RECT 9.7 0.45 10 1.95 ;
        RECT 0.6 0.45 0.9 10.95 ;
        RECT 4.9 9.45 8.8 9.75 ;
        RECT 8.5 8.85 8.8 9.75 ;
        RECT 1.8 4.05 2.7 4.35 ;
        RECT 1.8 1.05 2.1 4.95 ;
      LAYER Metal2 ;
        RECT 7.9 9.45 8.2 10.95 ;
        RECT 0.6 4.05 2.1 4.35 ;
      LAYER VIA1 ;
        RECT 0.65 4.1 0.85 4.3 ;
        RECT 1.85 4.1 2.05 4.3 ;
        RECT 7.95 10.7 8.15 10.9 ;
        RECT 7.95 9.5 8.15 9.7 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 18.5 0.15 ;
        RECT 1.2 10.05 17.9 10.35 ;
        RECT 17.6 -0.15 17.9 10.35 ;
        RECT 12.8 8.25 13.1 9.75 ;
        RECT 11.6 8.85 13.1 9.15 ;
        RECT 12.2 8.85 12.5 10.35 ;
        RECT 11.6 8.25 11.9 9.75 ;
        RECT 9.8 7.05 10.7 7.35 ;
        RECT 10.4 5.85 10.7 7.35 ;
        RECT 9.8 7.05 10.1 10.35 ;
        RECT 1.8 5.85 6.4 6.15 ;
        RECT 1.8 9.45 4 9.75 ;
        RECT 1.8 5.85 2.1 9.75 ;
        RECT 1.2 8.25 2.1 8.55 ;
        RECT 1.2 1.05 1.5 10.35 ;
        RECT 12.1 4.65 16.7 4.95 ;
        RECT 16.4 1.05 16.7 4.95 ;
        RECT 14.5 1.05 16.7 1.35 ;
        RECT 16.4 5.85 16.7 9.75 ;
        RECT 15.8 6.45 16.7 6.75 ;
        RECT 7.8 3.45 8.7 3.75 ;
        RECT 8.4 1.65 8.7 3.75 ;
        RECT 7.8 3.45 8.1 4.95 ;
        RECT 6.6 1.05 6.9 2.55 ;
        RECT 5.4 1.65 6.9 1.95 ;
        RECT 5.4 1.05 5.7 2.55 ;
      LAYER Metal2 ;
        RECT 16.4 1.05 17.9 1.35 ;
        RECT 16.4 6.45 17.9 6.75 ;
        RECT 8.4 -0.15 8.7 1.95 ;
        RECT 5.99 -0.15 6.29 1.95 ;
      LAYER VIA1 ;
        RECT 6.04 1.7 6.24 1.9 ;
        RECT 6.04 -0.1 6.24 0.1 ;
        RECT 8.45 1.7 8.65 1.9 ;
        RECT 8.45 -0.1 8.65 0.1 ;
        RECT 16.45 6.5 16.65 6.7 ;
        RECT 16.45 1.1 16.65 1.3 ;
        RECT 17.65 6.5 17.85 6.7 ;
        RECT 17.65 1.1 17.85 1.3 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 15.8 7.65 16.1 8.75 ;
      RECT 15.2 7.65 16.1 7.95 ;
      RECT 15.2 5.85 15.5 7.95 ;
      RECT 14 5.85 14.3 7.35 ;
      RECT 14 6.45 15.5 6.75 ;
      RECT 9.7 4.65 11.8 4.95 ;
      RECT 11.5 3.45 11.8 4.95 ;
      RECT 11.5 3.45 13.6 3.75 ;
      RECT 12.8 5.85 13.1 7.35 ;
      RECT 11.6 5.85 11.9 7.35 ;
      RECT 11.6 6.45 13.1 6.75 ;
      RECT 9.7 3.45 11.2 3.75 ;
      RECT 10.3 2.25 10.6 3.75 ;
      RECT 9.7 2.25 11.8 2.55 ;
      RECT 11.5 1.65 11.8 2.55 ;
      RECT 11.5 1.65 12.4 1.95 ;
      RECT 4.9 7.05 7 7.35 ;
      RECT 6.7 5.85 7 7.35 ;
      RECT 6.7 5.85 8.8 6.15 ;
      RECT 6.1 8.85 7 9.15 ;
      RECT 6.7 8.25 7 9.15 ;
      RECT 6.7 8.25 8.8 8.55 ;
      RECT 7.9 7.05 8.2 8.55 ;
      RECT 7.3 7.05 8.8 7.35 ;
      RECT 6.6 3.45 6.9 4.95 ;
      RECT 5.4 3.45 5.7 4.95 ;
      RECT 5.4 4.05 6.9 4.35 ;
      RECT 4.2 3.45 4.5 4.95 ;
      RECT 3 2.85 3.3 4.95 ;
      RECT 3 4.05 4.5 4.35 ;
      RECT 2.4 2.85 3.3 3.15 ;
      RECT 2.4 2.05 2.7 3.15 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END NAND2_1

MACRO NOR2_1
  CLASS CORE ;
  ORIGIN 0 0.15 ;
  FOREIGN NOR2_1 0 -0.15 ;
  SIZE 18.3 BY 11.1 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 12.6 1.65 14.1 1.95 ;
        RECT 13.2 5.85 13.5 7.35 ;
        RECT 4.2 8.85 5.7 9.15 ;
        RECT 4.8 3.45 5.1 4.95 ;
      LAYER Metal2 ;
        RECT 13.2 1.65 13.5 7.35 ;
        RECT 4.8 5.55 13.5 5.85 ;
        RECT 4.8 3.45 5.1 9.15 ;
      LAYER VIA1 ;
        RECT 4.85 8.9 5.05 9.1 ;
        RECT 4.85 4.1 5.05 4.3 ;
        RECT 13.25 6.5 13.45 6.7 ;
        RECT 13.25 1.7 13.45 1.9 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9 4.65 9.3 5.25 ;
      LAYER Metal2 ;
        RECT 8.7 4.95 12.9 5.25 ;
        RECT 12.6 4.35 12.9 5.25 ;
      LAYER VIA1 ;
        RECT 9.05 5 9.25 5.2 ;
    END
  END B
  PIN CTRL0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 6.6 7.65 6.9 7.95 ;
      LAYER Metal2 ;
        RECT 6.6 7.65 7.5 7.95 ;
        RECT 6.6 7.35 6.9 7.95 ;
      LAYER VIA1 ;
        RECT 6.65 7.7 6.85 7.9 ;
    END
  END CTRL0
  PIN CTRL1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 9.6 7.65 9.9 7.95 ;
      LAYER Metal2 ;
        RECT 9.6 7.65 10.5 7.95 ;
        RECT 9.6 7.05 9.9 7.95 ;
      LAYER VIA1 ;
        RECT 9.65 7.7 9.85 7.9 ;
    END
  END CTRL1
  PIN CTRL2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 15 2.85 15.3 3.15 ;
      LAYER Metal2 ;
        RECT 15 2.85 15.9 3.15 ;
        RECT 15 2.55 15.3 3.15 ;
      LAYER VIA1 ;
        RECT 15.05 2.9 15.25 3.1 ;
    END
  END CTRL2
  PIN CTRL3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 8.4 2.85 8.7 3.15 ;
      LAYER Metal2 ;
        RECT 8.1 2.85 8.7 3.15 ;
        RECT 8.4 2.25 8.7 3.15 ;
      LAYER VIA1 ;
        RECT 8.45 2.9 8.65 3.1 ;
    END
  END CTRL3
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal1 ;
        RECT 15 5.85 15.3 7.35 ;
        RECT 13.8 6.45 15.3 6.75 ;
        RECT 13.8 5.25 14.1 7.35 ;
        RECT 10.2 5.25 14.1 5.55 ;
        RECT 10.2 5.25 10.5 7.35 ;
        RECT 10.2 3.45 14.1 3.75 ;
        RECT 10.2 2.25 11.7 2.55 ;
        RECT 10.8 2.25 11.1 3.75 ;
        RECT 4.2 5.25 8.1 5.55 ;
        RECT 7.8 3.45 8.1 5.55 ;
        RECT 4.2 3.45 4.5 5.55 ;
        RECT 3 4.05 4.5 4.35 ;
        RECT 3 3.45 3.3 4.95 ;
        RECT 6.6 8.25 8.1 8.55 ;
        RECT 4.2 7.05 8.1 7.35 ;
        RECT 7.2 7.05 7.5 8.55 ;
      LAYER Metal2 ;
        RECT 3.6 9.45 14.7 9.75 ;
        RECT 14.4 3.45 14.7 9.75 ;
        RECT 13.8 3.45 14.7 3.75 ;
        RECT 3.6 7.05 4.5 7.35 ;
        RECT 3.6 4.05 3.9 9.75 ;
      LAYER VIA1 ;
        RECT 3.65 4.1 3.85 4.3 ;
        RECT 4.25 7.1 4.45 7.3 ;
        RECT 13.85 3.5 14.05 3.7 ;
        RECT 14.45 6.5 14.65 6.7 ;
    END
  END OUT
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 10.65 18.3 10.95 ;
        RECT 17.4 0.45 17.7 10.95 ;
        RECT 1.2 0.45 17.7 0.75 ;
        RECT 1.8 1.65 2.7 1.96 ;
        RECT 1.8 0.45 2.1 4.95 ;
        RECT 1.2 0.45 1.5 9.75 ;
        RECT 1.8 5.85 5.7 6.15 ;
        RECT 1.8 5.85 2.1 6.75 ;
      LAYER Metal2 ;
        RECT 1.2 5.85 2.3 6.15 ;
      LAYER VIA1 ;
        RECT 1.25 5.9 1.45 6.1 ;
        RECT 2.05 5.9 2.25 6.1 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal1 ;
        RECT 0 -0.15 18.3 0.15 ;
        RECT 0.6 10.05 17.1 10.35 ;
        RECT 16.8 1.05 17.1 10.35 ;
        RECT 12.6 4.65 17.1 4.95 ;
        RECT 16.2 5.85 16.5 10.35 ;
        RECT 16.2 4.05 16.5 4.95 ;
        RECT 15.6 8.84 16.5 9.15 ;
        RECT 12.6 8.25 12.9 9.75 ;
        RECT 11.4 8.85 12.9 9.15 ;
        RECT 12 8.85 12.3 10.35 ;
        RECT 11.4 8.25 11.7 9.75 ;
        RECT 1.8 9.45 8.7 9.75 ;
        RECT 8.4 5.85 8.7 9.75 ;
        RECT 6.6 5.85 8.7 6.15 ;
        RECT 4.8 9.45 5.1 10.35 ;
        RECT 0.6 -0.15 0.9 10.35 ;
        RECT 9.6 1.05 16.5 1.35 ;
        RECT 9.6 4.65 11.7 4.95 ;
        RECT 9.6 1.05 9.9 4.95 ;
        RECT 12.6 5.85 12.9 7.35 ;
        RECT 11.4 6.45 12.9 6.75 ;
        RECT 11.4 5.85 11.7 7.35 ;
        RECT 6.6 1.05 6.9 2.55 ;
        RECT 5.4 1.65 6.9 1.95 ;
        RECT 5.4 1.05 5.7 2.55 ;
        RECT 6.6 3.45 6.9 4.95 ;
        RECT 5.4 4.05 6.9 4.35 ;
        RECT 5.4 3.45 5.7 4.95 ;
      LAYER Metal2 ;
        RECT 15.6 -0.15 15.9 1.35 ;
        RECT 12 6.45 12.3 9.15 ;
        RECT 6 -0.15 6.3 4.35 ;
      LAYER VIA1 ;
        RECT 6.05 4.1 6.25 4.3 ;
        RECT 6.05 1.7 6.25 1.9 ;
        RECT 6.05 -0.1 6.25 0.1 ;
        RECT 12.05 8.9 12.25 9.1 ;
        RECT 12.05 6.5 12.25 6.7 ;
        RECT 15.65 1.1 15.85 1.3 ;
        RECT 15.65 -0.1 15.85 0.1 ;
    END
  END VSS
  OBS
    LAYER Metal1 ;
      RECT 13.8 4.05 14.7 4.35 ;
      RECT 14.4 3.45 14.7 4.35 ;
      RECT 14.4 3.45 16.5 3.75 ;
      RECT 15.6 2.25 15.9 3.75 ;
      RECT 12.6 2.25 16.5 2.55 ;
      RECT 15 7.65 15.3 9.75 ;
      RECT 13.8 7.65 14.1 9.75 ;
      RECT 10.2 7.65 10.5 9.75 ;
      RECT 13.8 8.85 15.3 9.15 ;
      RECT 15 7.65 15.9 7.95 ;
      RECT 15.6 6.85 15.9 7.95 ;
      RECT 10.2 7.65 14.1 7.95 ;
      RECT 2.4 2.85 2.7 3.95 ;
      RECT 4.2 2.85 8.1 3.15 ;
      RECT 7.8 1.05 8.1 3.15 ;
      RECT 2.4 2.85 3.3 3.15 ;
      RECT 3 1.05 3.3 3.15 ;
      RECT 4.2 1.05 4.5 3.15 ;
      RECT 3 1.65 4.5 1.95 ;
      RECT 1.8 8.25 5.7 8.55 ;
      RECT 2.4 7.05 2.7 8.55 ;
      RECT 1.8 7.05 3.9 7.35 ;
      RECT 3.6 6.45 3.9 7.35 ;
      RECT 3.6 6.45 4.5 6.75 ;
  END
  PROPERTY CatenaDesignType "deviceLevel" ;
END NOR2_1

END LIBRARY
